module multiply (output C,input A,input B);
assign C=A*B;
endmodule
