module multiply (output c,input a,input b);
assign c=a*b;
endmodule