package registr_param;
	parameter WIDTH_OUT                                  = 17;
endpackage