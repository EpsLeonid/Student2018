package V1_parameter;
parameter S=8;
endpackage
