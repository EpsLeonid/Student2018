package v4_param;

parameter k = 9;
parameter l = 5;
parameter M = 16;
parameter SIZE_IN = 17;
parameter SIZE_REG = 17;
parameter SIZE_OUT = 17;

endpackage
