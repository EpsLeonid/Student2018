package v2_parameter;
	parameter Vk = 5;
	parameter Vl = 5;
	parameter DELAY = Vk+Vl;
	parameter VM = 16;
endpackage