package parameters;
parameter N = 8;
endpackage 