package v2_parameter;
	parameter Vk = 5;
	parameter DELAY = k+1;
	parameter Vl = 5;
	parameter VM = 16;
endpackage