package v6_param;

parameter l = 6;
parameter k = 13;
parameter m1 = 16;
parameter m2 = 1;
parameter SIZE_IN = 17;
parameter SIZE_REG = 17;
parameter SIZE_OUT = 17;

endpackage
