package param_registr;

parameter WIDTH_OUT                                  = 17;

endpackage 