package parametr;
	parameter size = 8;
	parameter outsize = 16;

endpackage