package V2_param;

	parameter k = 5;
	parameter l = 5;
	parameter M = 16;
endpackage