package v5_parameter;

	parameter k                                     = 6;
	parameter l                                     = 6;
	parameter M                                     = 16;
	parameter DELAY                                 = k+l;

endpackage 