//---------------------
// ��������� ������� �1
// N=K+L

package v1_parameter;
parameter N_v1 =13;
parameter K_v1 =8;
parameter L_v1 =5;
parameter M_v1 =16;
endpackage