package v2_param;
	parameter V2_WIDTH= 16;
	parameter V2_k = 5;
	parameter V2_l = 5;
	parameter V2_M = 16;
endpackage