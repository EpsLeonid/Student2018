module verilog (
  input wire                   a,
  input wire                   b,
//--------------------------------
  output wire                  c);
//--------------------------------
  assign c=                   a&b;
//--------------------------------
endmodule
 