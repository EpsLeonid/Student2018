package parameters_v5;

parameter WIDTH_OUT                                  = 17;

endpackage 