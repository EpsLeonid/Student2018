package param;

	parameter WIDTH=17;
	
endpackage 