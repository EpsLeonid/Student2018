package v2_parameter;
	parameter Vk = 5;
	parameter DELAY = Vk+1;
	parameter Vl = 5;
	parameter VM = 16;
endpackage