package V2_param;
	parameter WIDTH = 16;
	parameter k = 5;
	parameter l = 5;
	parameter M = 16;
endpackage