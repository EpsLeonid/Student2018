module task1 (A, B, C);
	
	input wire A, B;
	output wire C;
	
	assign C = A * B;
endmodule 