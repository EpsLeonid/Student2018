package parameter;

	parameter WIDTH=17;
	
endpackage 