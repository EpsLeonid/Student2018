parameter WIDTH= 16;